module audio_lookback(
    input clk,                    
    input reset_n,  
    input button_s1,             // ��ťS1���� - δʹ��
    input button_s2,             // ��ťS2���� - δʹ��
    input button_s3,             // ��ťS3���� - ������С
    input button_s4,             // ��ťS4���� - ��������
    input uart_rx,               // ���ڽ���
    output reg led1,             // ��������ָʾ��LED1
    output reg led2,             // ����ָʾ��LED2
    output reg led3,             // ����Ч��ָʾ��LED3
    output reg led4,             // ��������ָʾ��LED4
    output reg led5,             // ������Сָʾ��LED5
    output led0,                 // ��ʼ�����ָʾ��LED0
                                  
    inout iic_0_scl,              
    inout iic_0_sda,   
    
    input I2S_DI,
    output I2S_RCLK,
    output I2S_BCLK,
    output I2S_DO,
    output I2S_MCLK
);

    parameter DATA_WIDTH = 32;     

    wire locked;
    
    // ʱ������
    clk_wiz_0 instance_name
    (
        .clk_out1(I2S_MCLK),     // output clk_out1
        .resetn(reset_n),        // input resetn
        .locked(locked),         // output locked
        .clk_in1(clk)            // input clk_in1
    );
    
    // BCLK��Ƶ
    clk_div4 clk_div4(
        .clk_in(I2S_MCLK),       // ����ʱ��
        .rst_n(reset_n),         // ��λ�ź�
        .clk_out(I2S_BCLK)       // ���ʱ��
    );

    // LRCK����
    reg[10:0] lrclk_cnt;
    reg i2s_lrck;
    always@(negedge I2S_BCLK or negedge reset_n)
    if(!reset_n) begin
        lrclk_cnt <= 11'd0;
        i2s_lrck <= 1'd0;
    end
    else if(~locked) begin
        lrclk_cnt <= 11'd0;
        i2s_lrck <= 1'd0;
    end
    else if(lrclk_cnt == 11'd64 - 1) begin          
        lrclk_cnt <= 11'd0;
        i2s_lrck <= ~i2s_lrck;
    end
    else begin
        lrclk_cnt <= lrclk_cnt + 1'd1;
        i2s_lrck <= i2s_lrck;
    end

    assign I2S_RCLK = i2s_lrck;

    // ES8388��ʼ��
    wire Init_Done;
    es8388_Init es8388_Init(
        .Clk(clk),
        .Rst_n(reset_n),
        .I2C_Init_Done(Init_Done),
        .i2c_sclk(iic_0_scl),
        .i2c_sdat(iic_0_sda)
    );
    
    assign led0 = Init_Done;

    // ���ڽ�������ź�
    wire [7:0] rx_data_byte;
    wire byte_rx_done;
    reg uart_echo_enable;        // ���ڿ��ƵĻ�������ʹ��
    reg uart_noise_reduction_enable; // ���ڿ��ƵĽ���ʹ��
    reg uart_echo_effect_enable;     // ���ڿ��ƵĻ���Ч��ʹ��
    
    // ����������������ź�
    reg uart_volume_up;
    reg uart_volume_down;
    reg [23:0] uart_volume_up_led_counter;
    reg [23:0] uart_volume_down_led_counter;
    reg uart_volume_up_led;
    reg uart_volume_down_led;
    
    // ���ڽ���ģ��ʵ����
    uart_byte_rx uart_rx_inst(
        .Clk(clk),
        .Rst_n(reset_n),
        .baud_set(3'd4),         // 115200������
        .uart_rx(uart_rx),
        .data_byte(rx_data_byte),
        .Rx_Done(byte_rx_done)
    );
    
    // ���������
    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            uart_echo_enable <= 1'b0;
            uart_noise_reduction_enable <= 1'b0;
            uart_echo_effect_enable <= 1'b0;
            uart_volume_up <= 1'b0;
            uart_volume_down <= 1'b0;
            uart_volume_up_led_counter <= 24'd0;
            uart_volume_down_led_counter <= 24'd0;
            uart_volume_up_led <= 1'b0;
            uart_volume_down_led <= 1'b0;
        end else begin
            // ��������LED������
            if (uart_volume_up_led_counter > 0) begin
                uart_volume_up_led_counter <= uart_volume_up_led_counter - 1'b1;
                uart_volume_up_led <= 1'b1;
            end else begin
                uart_volume_up_led <= 1'b0;
            end
            
            if (uart_volume_down_led_counter > 0) begin
                uart_volume_down_led_counter <= uart_volume_down_led_counter - 1'b1;
                uart_volume_down_led <= 1'b1;
            end else begin
                uart_volume_down_led <= 1'b0;
            end
            
            // ���������
            if (byte_rx_done) begin
                case(rx_data_byte)
                    8'h01: uart_echo_enable <= ~uart_echo_enable;           // �л���������״̬
                    8'h02: uart_noise_reduction_enable <= ~uart_noise_reduction_enable; // �л�����״̬
                    8'h03: uart_echo_effect_enable <= ~uart_echo_effect_enable;         // �л�����Ч��״̬
                    8'h0E: begin // 14 - ��������
                        uart_volume_up <= 1'b1;
                        uart_volume_up_led_counter <= 24'd2500000; // 50ms����
                    end
                    8'h0F: begin // 15 - ��С����
                        uart_volume_down <= 1'b1;
                        uart_volume_down_led_counter <= 24'd2500000; // 50ms����
                    end
                    default: begin
                        // �������������
                    end
                endcase
            end else begin
                // ����һ����������������������ź�
                uart_volume_up <= 1'b0;
                uart_volume_down <= 1'b0;
            end
        end
    end

    // ������������ź�
    wire volume_up_led;
    wire volume_down_led;
    wire [3:0] volume_level;     // 4λ֧��0-9����
    wire signed [15:0] volume_adjusted_left;
    wire signed [15:0] volume_adjusted_right;
    
    // ���յ�ʹ���źţ����ɴ��ڿ��ƣ�
    wire final_echo_enable = uart_echo_enable;
    wire final_noise_reduction_enable = uart_noise_reduction_enable;
    wire final_echo_effect_enable = uart_echo_effect_enable;
    
    // �ϲ�LEDָʾ�ź�
    wire combined_volume_up_led = volume_up_led | uart_volume_up_led;
    wire combined_volume_down_led = volume_down_led | uart_volume_down_led;
    
    // LED���ƺ�״̬�Ĵ���
    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            // LEDָʾ�Ƴ�ʼ��
            led1 <= 1'b0;
            led2 <= 1'b0;
            led3 <= 1'b0;
            led4 <= 1'b0;
            led5 <= 1'b0;
        end else begin
            // LED���ƣ����ɴ��ڿ���
            led1 <= final_echo_enable;           // LED1 - ��������
            led2 <= final_noise_reduction_enable; // LED2 - ����
            led3 <= final_echo_effect_enable;    // LED3 - ����Ч��
            
            // ��������LEDָʾ���ϲ���ť�ʹ��ڣ�
            led4 <= combined_volume_up_led;      // LED4 - ��������ָʾ
            led5 <= combined_volume_down_led;    // LED5 - ������Сָʾ
        end
    end

    // ��Ƶ���ݴ���
    reg adcfifo_read;
    wire [DATA_WIDTH - 1:0] adcfifo_readdata;
    wire adcfifo_empty;

    reg dacfifo_write;
    reg [DATA_WIDTH - 1:0] dacfifo_writedata;
    wire dacfifo_full;
    
    // ������������ź�
    wire signed [15:0] echo_data_out_left;
    wire signed [15:0] echo_data_out_right;
    
    // ��������ź�
    wire signed [15:0] noise_reduced_left;
    wire signed [15:0] noise_reduced_right;
    
    // �µĻ���Ч������ź�
    wire signed [15:0] echo_effect_left;
    wire signed [15:0] echo_effect_right;
    wire echo_effect_valid;
    
    // �м䴦���ź�
    wire signed [15:0] processed_left;
    wire signed [15:0] processed_right;
    
    // ��������ģ��ʵ����
    echo_cancellation echo_cancellation_inst (
        .sck(I2S_BCLK),
        .clk(clk),
        .rst_n(reset_n),
        .echo_enable(final_echo_enable),
        .data_in_left(adcfifo_readdata[31:16]),
        .data_in_right(adcfifo_readdata[15:0]),
        .data_out_left(echo_data_out_left),
        .data_out_right(echo_data_out_right)
    );
    
    // ѡ���������������ݻ�ԭʼ����
    assign processed_left = final_echo_enable ? echo_data_out_left : adcfifo_readdata[31:16];
    assign processed_right = final_echo_enable ? echo_data_out_right : adcfifo_readdata[15:0];
    
    // ����ģ��ʵ���� - ������
    advanced_noise_reduction noise_reduction_left (
        .clk(clk),
        .sck(I2S_BCLK),
        .rst_n(reset_n),
        .noise_reduction_enable(final_noise_reduction_enable),
        .data_in(processed_left),
        .data_out(noise_reduced_left)
    );
    
    // ����ģ��ʵ���� - ������
    advanced_noise_reduction noise_reduction_right (
        .clk(clk),
        .sck(I2S_BCLK),
        .rst_n(reset_n),
        .noise_reduction_enable(final_noise_reduction_enable),
        .data_in(processed_right),
        .data_out(noise_reduced_right)
    );
    
    // �������Ч��ģ��ʵ����
    simple_echo_effect echo_effect_inst (
        .clk(clk),
        .sck(I2S_BCLK),
        .rst_n(reset_n),
        .echo_effect_enable(final_echo_effect_enable),
        .data_in_left(noise_reduced_left),
        .data_in_right(noise_reduced_right),
        .data_valid(adcfifo_read),
        .data_out_left(echo_effect_left),
        .data_out_right(echo_effect_right),
        .data_out_valid(echo_effect_valid)
    );
        
    // ��������ģ��ʵ����
    volume_control volume_control_inst (
        .clk(clk),
        .sck(I2S_BCLK),
        .rst_n(reset_n),
        .volume_up(button_s4),           // S4������������
        .volume_down(button_s3),         // S3����������С
        .uart_volume_up(uart_volume_up), // ������������
        .uart_volume_down(uart_volume_down), // ����������С
        .data_in_left(final_echo_effect_enable ? echo_effect_left : noise_reduced_left),
        .data_in_right(final_echo_effect_enable ? echo_effect_right : noise_reduced_right),
        .data_out_left(volume_adjusted_left),
        .data_out_right(volume_adjusted_right),
        .volume_level(volume_level),
        .volume_up_led(volume_up_led),
        .volume_down_led(volume_down_led)
    );
    
    // ��������ѡ��
    always @(*) begin
        dacfifo_writedata = {volume_adjusted_left, volume_adjusted_right};
    end

    // ADC FIFO��ȡ����
    always @ (posedge clk or negedge reset_n)
    begin
        if (~reset_n)
        begin
            adcfifo_read <= 1'b0;
        end
        else if (~adcfifo_empty)
        begin
            adcfifo_read <= 1'b1;
        end
        else
        begin
            adcfifo_read <= 1'b0;
        end
    end

    // DAC FIFOд�����
    always @ (posedge clk or negedge reset_n)
    begin
        if(~reset_n)
            dacfifo_write <= 1'd0;
        else if(~dacfifo_full && (~adcfifo_empty)) begin
            dacfifo_write <= 1'd1;
        end
        else begin
            dacfifo_write <= 1'd0;
        end
    end

    // I2S����ģ��
    i2s_rx 
    #(
        .DATA_WIDTH(DATA_WIDTH) 
    ) i2s_rx_inst
    (
        .reset_n(reset_n),
        .bclk(I2S_BCLK),
        .adclrc(I2S_RCLK),
        .adcdat(I2S_DI),
        .adcfifo_rdclk(clk),
        .adcfifo_read(adcfifo_read),
        .adcfifo_empty(adcfifo_empty),
        .adcfifo_readdata(adcfifo_readdata)
    );
    
    // I2S����ģ��
    i2s_tx
    #(
         .DATA_WIDTH(DATA_WIDTH)
    ) i2s_tx_inst
    (
         .reset_n(reset_n),
         .dacfifo_wrclk(clk),
         .dacfifo_wren(dacfifo_write),
         .dacfifo_wrdata(dacfifo_writedata),
         .dacfifo_full(dacfifo_full),
         .bclk(I2S_BCLK),
         .daclrc(I2S_RCLK),
         .dacdat(I2S_DO)
    );

endmodule